module tb_decoder_4line_16line();
	reg [3:0] sel;
	wire [15:0] out;
endmodule
