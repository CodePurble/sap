module main();
endmodule
